// vga_lt24_accelerometer_computer.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module vga_lt24_accelerometer_computer (
		inout  wire        accelerometer_spi_export_I2C_SDAT,          //            accelerometer_spi_export.I2C_SDAT
		output wire        accelerometer_spi_export_I2C_SCLK,          //                                    .I2C_SCLK
		output wire        accelerometer_spi_export_G_SENSOR_CS_N,     //                                    .G_SENSOR_CS_N
		input  wire        accelerometer_spi_export_G_SENSOR_INT,      //                                    .G_SENSOR_INT
		input  wire        clk_clk,                                    //                                 clk.clk
		output wire [31:0] hex3_hex0_out_export,                       //                       hex3_hex0_out.export
		output wire [15:0] hex5_hex4_out_export,                       //                       hex5_hex4_out.export
		input  wire [1:0]  key_out_export,                             //                             key_out.export
		output wire        lcd_reset_n_external_connection_export,     //     lcd_reset_n_external_connection.export
		output wire [9:0]  leds_out_export,                            //                            leds_out.export
		output wire        lt24_controller_conduit_end_cs,             //         lt24_controller_conduit_end.cs
		output wire        lt24_controller_conduit_end_rs,             //                                    .rs
		output wire        lt24_controller_conduit_end_rd,             //                                    .rd
		output wire        lt24_controller_conduit_end_wr,             //                                    .wr
		output wire [15:0] lt24_controller_conduit_end_data,           //                                    .data
		input  wire        reset_reset_n,                              //                               reset.reset_n
		output wire        sdram_clk_clk,                              //                           sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                            //                          sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                              //                                    .ba
		output wire        sdram_wire_cas_n,                           //                                    .cas_n
		output wire        sdram_wire_cke,                             //                                    .cke
		output wire        sdram_wire_cs_n,                            //                                    .cs_n
		inout  wire [15:0] sdram_wire_dq,                              //                                    .dq
		output wire [1:0]  sdram_wire_dqm,                             //                                    .dqm
		output wire        sdram_wire_ras_n,                           //                                    .ras_n
		output wire        sdram_wire_we_n,                            //                                    .we_n
		input  wire [9:0]  sliders_out_export,                         //                         sliders_out.export
		input  wire        spi_external_MISO,                          //                        spi_external.MISO
		output wire        spi_external_MOSI,                          //                                    .MOSI
		output wire        spi_external_SCLK,                          //                                    .SCLK
		output wire        spi_external_SS_n,                          //                                    .SS_n
		input  wire        touch_busy_external_connection_export,      //      touch_busy_external_connection.export
		input  wire        touch_pen_irq_n_external_connection_export, // touch_pen_irq_n_external_connection.export
		output wire        vga_output_CLK,                             //                          vga_output.CLK
		output wire        vga_output_HS,                              //                                    .HS
		output wire        vga_output_VS,                              //                                    .VS
		output wire        vga_output_BLANK,                           //                                    .BLANK
		output wire        vga_output_SYNC,                            //                                    .SYNC
		output wire [3:0]  vga_output_R,                               //                                    .R
		output wire [3:0]  vga_output_G,                               //                                    .G
		output wire [3:0]  vga_output_B                                //                                    .B
	);

	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_valid;                             // video_dual_clock_buffer_0:stream_out_valid -> video_vga_controller_0:valid
	wire  [29:0] video_dual_clock_buffer_0_avalon_dc_buffer_source_data;                              // video_dual_clock_buffer_0:stream_out_data -> video_vga_controller_0:data
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_ready;                             // video_vga_controller_0:ready -> video_dual_clock_buffer_0:stream_out_ready
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket;                     // video_dual_clock_buffer_0:stream_out_startofpacket -> video_vga_controller_0:startofpacket
	wire         video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket;                       // video_dual_clock_buffer_0:stream_out_endofpacket -> video_vga_controller_0:endofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_valid;                                  // video_pixel_buffer_dma_0:stream_valid -> video_rgb_resampler_0:stream_in_valid
	wire  [15:0] video_pixel_buffer_dma_0_avalon_pixel_source_data;                                   // video_pixel_buffer_dma_0:stream_data -> video_rgb_resampler_0:stream_in_data
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_ready;                                  // video_rgb_resampler_0:stream_in_ready -> video_pixel_buffer_dma_0:stream_ready
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket;                          // video_pixel_buffer_dma_0:stream_startofpacket -> video_rgb_resampler_0:stream_in_startofpacket
	wire         video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket;                            // video_pixel_buffer_dma_0:stream_endofpacket -> video_rgb_resampler_0:stream_in_endofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_valid;                                       // video_rgb_resampler_0:stream_out_valid -> video_dual_clock_buffer_0:stream_in_valid
	wire  [29:0] video_rgb_resampler_0_avalon_rgb_source_data;                                        // video_rgb_resampler_0:stream_out_data -> video_dual_clock_buffer_0:stream_in_data
	wire         video_rgb_resampler_0_avalon_rgb_source_ready;                                       // video_dual_clock_buffer_0:stream_in_ready -> video_rgb_resampler_0:stream_out_ready
	wire         video_rgb_resampler_0_avalon_rgb_source_startofpacket;                               // video_rgb_resampler_0:stream_out_startofpacket -> video_dual_clock_buffer_0:stream_in_startofpacket
	wire         video_rgb_resampler_0_avalon_rgb_source_endofpacket;                                 // video_rgb_resampler_0:stream_out_endofpacket -> video_dual_clock_buffer_0:stream_in_endofpacket
	wire         altpll_0_c0_clk;                                                                     // altpll_0:c0 -> [rst_controller_004:clk, video_dual_clock_buffer_0:clk_stream_out, video_vga_controller_0:clk]
	wire         altpll_0_c2_clk;                                                                     // altpll_0:c2 -> [HEX3_HEX0:clk, HEX5_HEX4:clk, KEY:clk, LEDS:clk, LT24_Controller:clk, SLIDERS:clk, accelerometer_spi:clk, irq_mapper:clk, irq_synchronizer:sender_clk, irq_synchronizer_001:sender_clk, jtag_uart_0:clk, mm_clock_crossing_bridge:s0_clk, mm_interconnect_0:altpll_0_c2_clk, mm_interconnect_1:altpll_0_c2_clk, new_sdram_controller_0:clk, nios2_gen2_0:clk, onchip_memory2_0:clk, rst_controller:clk, rst_controller_002:clk, sysid_qsys_0:clock, timer_0:clk, timer_1:clk, video_dual_clock_buffer_0:clk_stream_in, video_pixel_buffer_dma_0:clk, video_rgb_resampler_0:clk]
	wire         altpll_0_c3_clk;                                                                     // altpll_0:c3 -> [LCD_RESET_N:clk, irq_synchronizer:receiver_clk, irq_synchronizer_001:receiver_clk, mm_clock_crossing_bridge:m0_clk, mm_interconnect_1:altpll_0_c3_clk, rst_controller_001:clk, touch_busy:clk, touch_pen_irq_n:clk, touch_spi:clk]
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest;                        // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest -> video_pixel_buffer_dma_0:master_waitrequest
	wire  [15:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata;                           // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata -> video_pixel_buffer_dma_0:master_readdata
	wire  [31:0] video_pixel_buffer_dma_0_avalon_pixel_dma_master_address;                            // video_pixel_buffer_dma_0:master_address -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_address
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_read;                               // video_pixel_buffer_dma_0:master_read -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_read
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid;                      // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid -> video_pixel_buffer_dma_0:master_readdatavalid
	wire         video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock;                               // video_pixel_buffer_dma_0:master_arbiterlock -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock
	wire  [31:0] nios2_gen2_0_data_master_readdata;                                                   // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                                                // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                                                // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [26:0] nios2_gen2_0_data_master_address;                                                    // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                                                 // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                                                       // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_readdatavalid;                                              // mm_interconnect_0:nios2_gen2_0_data_master_readdatavalid -> nios2_gen2_0:d_readdatavalid
	wire         nios2_gen2_0_data_master_write;                                                      // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                                                  // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire   [3:0] nios2_gen2_0_data_master_burstcount;                                                 // nios2_gen2_0:d_burstcount -> mm_interconnect_0:nios2_gen2_0_data_master_burstcount
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                                            // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                                         // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [26:0] nios2_gen2_0_instruction_master_address;                                             // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                                                // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         nios2_gen2_0_instruction_master_readdatavalid;                                       // mm_interconnect_0:nios2_gen2_0_instruction_master_readdatavalid -> nios2_gen2_0:i_readdatavalid
	wire   [3:0] nios2_gen2_0_instruction_master_burstcount;                                          // nios2_gen2_0:i_burstcount -> mm_interconnect_0:nios2_gen2_0_instruction_master_burstcount
	wire         mm_interconnect_0_new_sdram_controller_0_s1_chipselect;                              // mm_interconnect_0:new_sdram_controller_0_s1_chipselect -> new_sdram_controller_0:az_cs
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_readdata;                                // new_sdram_controller_0:za_data -> mm_interconnect_0:new_sdram_controller_0_s1_readdata
	wire         mm_interconnect_0_new_sdram_controller_0_s1_waitrequest;                             // new_sdram_controller_0:za_waitrequest -> mm_interconnect_0:new_sdram_controller_0_s1_waitrequest
	wire  [24:0] mm_interconnect_0_new_sdram_controller_0_s1_address;                                 // mm_interconnect_0:new_sdram_controller_0_s1_address -> new_sdram_controller_0:az_addr
	wire         mm_interconnect_0_new_sdram_controller_0_s1_read;                                    // mm_interconnect_0:new_sdram_controller_0_s1_read -> new_sdram_controller_0:az_rd_n
	wire   [1:0] mm_interconnect_0_new_sdram_controller_0_s1_byteenable;                              // mm_interconnect_0:new_sdram_controller_0_s1_byteenable -> new_sdram_controller_0:az_be_n
	wire         mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid;                           // new_sdram_controller_0:za_valid -> mm_interconnect_0:new_sdram_controller_0_s1_readdatavalid
	wire         mm_interconnect_0_new_sdram_controller_0_s1_write;                                   // mm_interconnect_0:new_sdram_controller_0_s1_write -> new_sdram_controller_0:az_wr_n
	wire  [15:0] mm_interconnect_0_new_sdram_controller_0_s1_writedata;                               // mm_interconnect_0:new_sdram_controller_0_s1_writedata -> new_sdram_controller_0:az_data
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;                             // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;                          // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;                          // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;                              // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;                                 // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;                           // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;                                // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;                            // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_chipselect;                                    // mm_interconnect_0:onchip_memory2_0_s1_chipselect -> onchip_memory2_0:chipselect
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_readdata;                                      // onchip_memory2_0:readdata -> mm_interconnect_0:onchip_memory2_0_s1_readdata
	wire   [7:0] mm_interconnect_0_onchip_memory2_0_s1_address;                                       // mm_interconnect_0:onchip_memory2_0_s1_address -> onchip_memory2_0:address
	wire   [3:0] mm_interconnect_0_onchip_memory2_0_s1_byteenable;                                    // mm_interconnect_0:onchip_memory2_0_s1_byteenable -> onchip_memory2_0:byteenable
	wire         mm_interconnect_0_onchip_memory2_0_s1_write;                                         // mm_interconnect_0:onchip_memory2_0_s1_write -> onchip_memory2_0:write
	wire  [31:0] mm_interconnect_0_onchip_memory2_0_s1_writedata;                                     // mm_interconnect_0:onchip_memory2_0_s1_writedata -> onchip_memory2_0:writedata
	wire         mm_interconnect_0_onchip_memory2_0_s1_clken;                                         // mm_interconnect_0:onchip_memory2_0_s1_clken -> onchip_memory2_0:clken
	wire   [7:0] mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_readdata;    // accelerometer_spi:readdata -> mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_readdata
	wire         mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_waitrequest; // accelerometer_spi:waitrequest -> mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_waitrequest
	wire   [0:0] mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_address;     // mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_address -> accelerometer_spi:address
	wire         mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_read;        // mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_read -> accelerometer_spi:read
	wire   [0:0] mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_byteenable;  // mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_byteenable -> accelerometer_spi:byteenable
	wire         mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_write;       // mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_write -> accelerometer_spi:write
	wire   [7:0] mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_writedata;   // mm_interconnect_0:accelerometer_spi_avalon_accelerometer_spi_mode_slave_writedata -> accelerometer_spi:writedata
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata;            // video_pixel_buffer_dma_0:slave_readdata -> mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_readdata
	wire   [1:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address;             // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_address -> video_pixel_buffer_dma_0:slave_address
	wire         mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read;                // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_read -> video_pixel_buffer_dma_0:slave_read
	wire   [3:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable;          // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_byteenable -> video_pixel_buffer_dma_0:slave_byteenable
	wire         mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write;               // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_write -> video_pixel_buffer_dma_0:slave_write
	wire  [31:0] mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata;           // mm_interconnect_0:video_pixel_buffer_dma_0_avalon_control_slave_writedata -> video_pixel_buffer_dma_0:slave_writedata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;                          // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;                            // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest;                         // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;                             // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;                                // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;                               // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;                           // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata;                   // video_rgb_resampler_0:slave_readdata -> mm_interconnect_0:video_rgb_resampler_0_avalon_rgb_slave_readdata
	wire         mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read;                       // mm_interconnect_0:video_rgb_resampler_0_avalon_rgb_slave_read -> video_rgb_resampler_0:slave_read
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;                               // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;                                // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;                                       // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;                                        // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                                           // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                                          // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;                                      // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata;                              // mm_clock_crossing_bridge:s0_readdata -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdata
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest;                           // mm_clock_crossing_bridge:s0_waitrequest -> mm_interconnect_0:mm_clock_crossing_bridge_s0_waitrequest
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess;                           // mm_interconnect_0:mm_clock_crossing_bridge_s0_debugaccess -> mm_clock_crossing_bridge:s0_debugaccess
	wire   [9:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_address;                               // mm_interconnect_0:mm_clock_crossing_bridge_s0_address -> mm_clock_crossing_bridge:s0_address
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_read;                                  // mm_interconnect_0:mm_clock_crossing_bridge_s0_read -> mm_clock_crossing_bridge:s0_read
	wire   [3:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable;                            // mm_interconnect_0:mm_clock_crossing_bridge_s0_byteenable -> mm_clock_crossing_bridge:s0_byteenable
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid;                         // mm_clock_crossing_bridge:s0_readdatavalid -> mm_interconnect_0:mm_clock_crossing_bridge_s0_readdatavalid
	wire         mm_interconnect_0_mm_clock_crossing_bridge_s0_write;                                 // mm_interconnect_0:mm_clock_crossing_bridge_s0_write -> mm_clock_crossing_bridge:s0_write
	wire  [31:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata;                             // mm_interconnect_0:mm_clock_crossing_bridge_s0_writedata -> mm_clock_crossing_bridge:s0_writedata
	wire   [0:0] mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount;                            // mm_interconnect_0:mm_clock_crossing_bridge_s0_burstcount -> mm_clock_crossing_bridge:s0_burstcount
	wire         mm_interconnect_0_timer_0_s1_chipselect;                                             // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                                               // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                                                // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                                                  // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                                              // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_key_s1_chipselect;                                                 // mm_interconnect_0:KEY_s1_chipselect -> KEY:chipselect
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                                                   // KEY:readdata -> mm_interconnect_0:KEY_s1_readdata
	wire   [1:0] mm_interconnect_0_key_s1_address;                                                    // mm_interconnect_0:KEY_s1_address -> KEY:address
	wire         mm_interconnect_0_key_s1_write;                                                      // mm_interconnect_0:KEY_s1_write -> KEY:write_n
	wire  [31:0] mm_interconnect_0_key_s1_writedata;                                                  // mm_interconnect_0:KEY_s1_writedata -> KEY:writedata
	wire  [31:0] mm_interconnect_0_sliders_s1_readdata;                                               // SLIDERS:readdata -> mm_interconnect_0:SLIDERS_s1_readdata
	wire   [1:0] mm_interconnect_0_sliders_s1_address;                                                // mm_interconnect_0:SLIDERS_s1_address -> SLIDERS:address
	wire         mm_interconnect_0_hex3_hex0_s1_chipselect;                                           // mm_interconnect_0:HEX3_HEX0_s1_chipselect -> HEX3_HEX0:chipselect
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_readdata;                                             // HEX3_HEX0:readdata -> mm_interconnect_0:HEX3_HEX0_s1_readdata
	wire   [1:0] mm_interconnect_0_hex3_hex0_s1_address;                                              // mm_interconnect_0:HEX3_HEX0_s1_address -> HEX3_HEX0:address
	wire         mm_interconnect_0_hex3_hex0_s1_write;                                                // mm_interconnect_0:HEX3_HEX0_s1_write -> HEX3_HEX0:write_n
	wire  [31:0] mm_interconnect_0_hex3_hex0_s1_writedata;                                            // mm_interconnect_0:HEX3_HEX0_s1_writedata -> HEX3_HEX0:writedata
	wire         mm_interconnect_0_hex5_hex4_s1_chipselect;                                           // mm_interconnect_0:HEX5_HEX4_s1_chipselect -> HEX5_HEX4:chipselect
	wire  [31:0] mm_interconnect_0_hex5_hex4_s1_readdata;                                             // HEX5_HEX4:readdata -> mm_interconnect_0:HEX5_HEX4_s1_readdata
	wire   [1:0] mm_interconnect_0_hex5_hex4_s1_address;                                              // mm_interconnect_0:HEX5_HEX4_s1_address -> HEX5_HEX4:address
	wire         mm_interconnect_0_hex5_hex4_s1_write;                                                // mm_interconnect_0:HEX5_HEX4_s1_write -> HEX5_HEX4:write_n
	wire  [31:0] mm_interconnect_0_hex5_hex4_s1_writedata;                                            // mm_interconnect_0:HEX5_HEX4_s1_writedata -> HEX5_HEX4:writedata
	wire         mm_interconnect_0_leds_s1_chipselect;                                                // mm_interconnect_0:LEDS_s1_chipselect -> LEDS:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                                                  // LEDS:readdata -> mm_interconnect_0:LEDS_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                                                   // mm_interconnect_0:LEDS_s1_address -> LEDS:address
	wire         mm_interconnect_0_leds_s1_write;                                                     // mm_interconnect_0:LEDS_s1_write -> LEDS:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                                                 // mm_interconnect_0:LEDS_s1_writedata -> LEDS:writedata
	wire         mm_interconnect_0_timer_1_s1_chipselect;                                             // mm_interconnect_0:timer_1_s1_chipselect -> timer_1:chipselect
	wire  [15:0] mm_interconnect_0_timer_1_s1_readdata;                                               // timer_1:readdata -> mm_interconnect_0:timer_1_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_1_s1_address;                                                // mm_interconnect_0:timer_1_s1_address -> timer_1:address
	wire         mm_interconnect_0_timer_1_s1_write;                                                  // mm_interconnect_0:timer_1_s1_write -> timer_1:write_n
	wire  [15:0] mm_interconnect_0_timer_1_s1_writedata;                                              // mm_interconnect_0:timer_1_s1_writedata -> timer_1:writedata
	wire         mm_clock_crossing_bridge_m0_waitrequest;                                             // mm_interconnect_1:mm_clock_crossing_bridge_m0_waitrequest -> mm_clock_crossing_bridge:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_m0_readdata;                                                // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdata -> mm_clock_crossing_bridge:m0_readdata
	wire         mm_clock_crossing_bridge_m0_debugaccess;                                             // mm_clock_crossing_bridge:m0_debugaccess -> mm_interconnect_1:mm_clock_crossing_bridge_m0_debugaccess
	wire   [9:0] mm_clock_crossing_bridge_m0_address;                                                 // mm_clock_crossing_bridge:m0_address -> mm_interconnect_1:mm_clock_crossing_bridge_m0_address
	wire         mm_clock_crossing_bridge_m0_read;                                                    // mm_clock_crossing_bridge:m0_read -> mm_interconnect_1:mm_clock_crossing_bridge_m0_read
	wire   [3:0] mm_clock_crossing_bridge_m0_byteenable;                                              // mm_clock_crossing_bridge:m0_byteenable -> mm_interconnect_1:mm_clock_crossing_bridge_m0_byteenable
	wire         mm_clock_crossing_bridge_m0_readdatavalid;                                           // mm_interconnect_1:mm_clock_crossing_bridge_m0_readdatavalid -> mm_clock_crossing_bridge:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_m0_writedata;                                               // mm_clock_crossing_bridge:m0_writedata -> mm_interconnect_1:mm_clock_crossing_bridge_m0_writedata
	wire         mm_clock_crossing_bridge_m0_write;                                                   // mm_clock_crossing_bridge:m0_write -> mm_interconnect_1:mm_clock_crossing_bridge_m0_write
	wire   [0:0] mm_clock_crossing_bridge_m0_burstcount;                                              // mm_clock_crossing_bridge:m0_burstcount -> mm_interconnect_1:mm_clock_crossing_bridge_m0_burstcount
	wire         mm_interconnect_1_lt24_controller_avalon_slave_0_chipselect;                         // mm_interconnect_1:LT24_Controller_avalon_slave_0_chipselect -> LT24_Controller:s_chipselect_n
	wire   [0:0] mm_interconnect_1_lt24_controller_avalon_slave_0_address;                            // mm_interconnect_1:LT24_Controller_avalon_slave_0_address -> LT24_Controller:s_address
	wire         mm_interconnect_1_lt24_controller_avalon_slave_0_write;                              // mm_interconnect_1:LT24_Controller_avalon_slave_0_write -> LT24_Controller:s_write_n
	wire  [31:0] mm_interconnect_1_lt24_controller_avalon_slave_0_writedata;                          // mm_interconnect_1:LT24_Controller_avalon_slave_0_writedata -> LT24_Controller:s_writedata
	wire         mm_interconnect_1_lcd_reset_n_s1_chipselect;                                         // mm_interconnect_1:LCD_RESET_N_s1_chipselect -> LCD_RESET_N:chipselect
	wire  [31:0] mm_interconnect_1_lcd_reset_n_s1_readdata;                                           // LCD_RESET_N:readdata -> mm_interconnect_1:LCD_RESET_N_s1_readdata
	wire   [1:0] mm_interconnect_1_lcd_reset_n_s1_address;                                            // mm_interconnect_1:LCD_RESET_N_s1_address -> LCD_RESET_N:address
	wire         mm_interconnect_1_lcd_reset_n_s1_write;                                              // mm_interconnect_1:LCD_RESET_N_s1_write -> LCD_RESET_N:write_n
	wire  [31:0] mm_interconnect_1_lcd_reset_n_s1_writedata;                                          // mm_interconnect_1:LCD_RESET_N_s1_writedata -> LCD_RESET_N:writedata
	wire         mm_interconnect_1_touch_pen_irq_n_s1_chipselect;                                     // mm_interconnect_1:touch_pen_irq_n_s1_chipselect -> touch_pen_irq_n:chipselect
	wire  [31:0] mm_interconnect_1_touch_pen_irq_n_s1_readdata;                                       // touch_pen_irq_n:readdata -> mm_interconnect_1:touch_pen_irq_n_s1_readdata
	wire   [1:0] mm_interconnect_1_touch_pen_irq_n_s1_address;                                        // mm_interconnect_1:touch_pen_irq_n_s1_address -> touch_pen_irq_n:address
	wire         mm_interconnect_1_touch_pen_irq_n_s1_write;                                          // mm_interconnect_1:touch_pen_irq_n_s1_write -> touch_pen_irq_n:write_n
	wire  [31:0] mm_interconnect_1_touch_pen_irq_n_s1_writedata;                                      // mm_interconnect_1:touch_pen_irq_n_s1_writedata -> touch_pen_irq_n:writedata
	wire  [31:0] mm_interconnect_1_touch_busy_s1_readdata;                                            // touch_busy:readdata -> mm_interconnect_1:touch_busy_s1_readdata
	wire   [1:0] mm_interconnect_1_touch_busy_s1_address;                                             // mm_interconnect_1:touch_busy_s1_address -> touch_busy:address
	wire         mm_interconnect_1_touch_spi_spi_control_port_chipselect;                             // mm_interconnect_1:touch_spi_spi_control_port_chipselect -> touch_spi:spi_select
	wire  [15:0] mm_interconnect_1_touch_spi_spi_control_port_readdata;                               // touch_spi:data_to_cpu -> mm_interconnect_1:touch_spi_spi_control_port_readdata
	wire   [2:0] mm_interconnect_1_touch_spi_spi_control_port_address;                                // mm_interconnect_1:touch_spi_spi_control_port_address -> touch_spi:mem_addr
	wire         mm_interconnect_1_touch_spi_spi_control_port_read;                                   // mm_interconnect_1:touch_spi_spi_control_port_read -> touch_spi:read_n
	wire         mm_interconnect_1_touch_spi_spi_control_port_write;                                  // mm_interconnect_1:touch_spi_spi_control_port_write -> touch_spi:write_n
	wire  [15:0] mm_interconnect_1_touch_spi_spi_control_port_writedata;                              // mm_interconnect_1:touch_spi_spi_control_port_writedata -> touch_spi:data_from_cpu
	wire         irq_mapper_receiver0_irq;                                                            // accelerometer_spi:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                            // jtag_uart_0:av_irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                            // timer_0:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver5_irq;                                                            // timer_1:irq -> irq_mapper:receiver5_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                                                // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         irq_mapper_receiver3_irq;                                                            // irq_synchronizer:sender_irq -> irq_mapper:receiver3_irq
	wire   [0:0] irq_synchronizer_receiver_irq;                                                       // touch_pen_irq_n:irq -> irq_synchronizer:receiver_irq
	wire         irq_mapper_receiver4_irq;                                                            // irq_synchronizer_001:sender_irq -> irq_mapper:receiver4_irq
	wire   [0:0] irq_synchronizer_001_receiver_irq;                                                   // touch_spi:irq -> irq_synchronizer_001:receiver_irq
	wire         rst_controller_reset_out_reset;                                                      // rst_controller:reset_out -> [HEX3_HEX0:reset_n, HEX5_HEX4:reset_n, KEY:reset_n, LEDS:reset_n, SLIDERS:reset_n, accelerometer_spi:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, jtag_uart_0:rst_n, mm_interconnect_0:video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset, new_sdram_controller_0:reset_n, nios2_gen2_0:reset_n, onchip_memory2_0:reset, rst_translator:in_reset, sysid_qsys_0:reset_n, timer_0:reset_n, video_dual_clock_buffer_0:reset_stream_in, video_pixel_buffer_dma_0:reset, video_rgb_resampler_0:reset]
	wire         rst_controller_reset_out_reset_req;                                                  // rst_controller:reset_req -> [nios2_gen2_0:reset_req, onchip_memory2_0:reset_req, rst_translator:reset_req_in]
	wire         nios2_gen2_0_debug_reset_request_reset;                                              // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_003:reset_in1, rst_controller_004:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                                  // rst_controller_001:reset_out -> [LCD_RESET_N:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, mm_clock_crossing_bridge:m0_reset, mm_interconnect_1:mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset, touch_busy:reset_n, touch_pen_irq_n:reset_n, touch_spi:reset_n]
	wire         rst_controller_002_reset_out_reset;                                                  // rst_controller_002:reset_out -> [LT24_Controller:reset_n, mm_clock_crossing_bridge:s0_reset, mm_interconnect_0:mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset_reset, mm_interconnect_1:LT24_Controller_reset_reset_bridge_in_reset_reset, timer_1:reset_n]
	wire         rst_controller_003_reset_out_reset;                                                  // rst_controller_003:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire         rst_controller_004_reset_out_reset;                                                  // rst_controller_004:reset_out -> [video_dual_clock_buffer_0:reset_stream_out, video_vga_controller_0:reset]

	vga_lt24_accelerometer_computer_HEX3_HEX0 hex3_hex0 (
		.clk        (altpll_0_c2_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex3_hex0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex3_hex0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex3_hex0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex3_hex0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex3_hex0_s1_readdata),   //                    .readdata
		.out_port   (hex3_hex0_out_export)                       // external_connection.export
	);

	vga_lt24_accelerometer_computer_HEX5_HEX4 hex5_hex4 (
		.clk        (altpll_0_c2_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_hex5_hex4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_hex5_hex4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_hex5_hex4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_hex5_hex4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_hex5_hex4_s1_readdata),   //                    .readdata
		.out_port   (hex5_hex4_out_export)                       // external_connection.export
	);

	vga_lt24_accelerometer_computer_KEY key (
		.clk        (altpll_0_c2_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (key_out_export)                       // external_connection.export
	);

	vga_lt24_accelerometer_computer_LCD_RESET_N lcd_reset_n (
		.clk        (altpll_0_c3_clk),                             //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_1_lcd_reset_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_lcd_reset_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_lcd_reset_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_lcd_reset_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_lcd_reset_n_s1_readdata),   //                    .readdata
		.out_port   (lcd_reset_n_external_connection_export)       // external_connection.export
	);

	vga_lt24_accelerometer_computer_LEDS leds (
		.clk        (altpll_0_c2_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_out_export)                       // external_connection.export
	);

	LT24_Controller lt24_controller (
		.clk            (altpll_0_c2_clk),                                              //          clock.clk
		.reset_n        (~rst_controller_002_reset_out_reset),                          //          reset.reset_n
		.s_chipselect_n (~mm_interconnect_1_lt24_controller_avalon_slave_0_chipselect), // avalon_slave_0.chipselect_n
		.s_write_n      (~mm_interconnect_1_lt24_controller_avalon_slave_0_write),      //               .write_n
		.s_writedata    (mm_interconnect_1_lt24_controller_avalon_slave_0_writedata),   //               .writedata
		.s_address      (mm_interconnect_1_lt24_controller_avalon_slave_0_address),     //               .address
		.lt24_cs        (lt24_controller_conduit_end_cs),                               //    conduit_end.export
		.lt24_rs        (lt24_controller_conduit_end_rs),                               //               .export
		.lt24_rd        (lt24_controller_conduit_end_rd),                               //               .export
		.lt24_wr        (lt24_controller_conduit_end_wr),                               //               .export
		.lt24_data      (lt24_controller_conduit_end_data)                              //               .export
	);

	vga_lt24_accelerometer_computer_SLIDERS sliders (
		.clk      (altpll_0_c2_clk),                       //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_sliders_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sliders_s1_readdata), //                    .readdata
		.in_port  (sliders_out_export)                     // external_connection.export
	);

	vga_lt24_accelerometer_computer_accelerometer_spi accelerometer_spi (
		.clk           (altpll_0_c2_clk),                                                                     //                                 clk.clk
		.reset         (rst_controller_reset_out_reset),                                                      //                               reset.reset
		.address       (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_address),     // avalon_accelerometer_spi_mode_slave.address
		.byteenable    (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_byteenable),  //                                    .byteenable
		.read          (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_read),        //                                    .read
		.write         (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_write),       //                                    .write
		.writedata     (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_writedata),   //                                    .writedata
		.readdata      (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_readdata),    //                                    .readdata
		.waitrequest   (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_waitrequest), //                                    .waitrequest
		.irq           (irq_mapper_receiver0_irq),                                                            //                           interrupt.irq
		.I2C_SDAT      (accelerometer_spi_export_I2C_SDAT),                                                   //                  external_interface.export
		.I2C_SCLK      (accelerometer_spi_export_I2C_SCLK),                                                   //                                    .export
		.G_SENSOR_CS_N (accelerometer_spi_export_G_SENSOR_CS_N),                                              //                                    .export
		.G_SENSOR_INT  (accelerometer_spi_export_G_SENSOR_INT)                                                //                                    .export
	);

	vga_lt24_accelerometer_computer_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_003_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                                  //                    c1.clk
		.c2                 (altpll_0_c2_clk),                                //                    c2.clk
		.c3                 (altpll_0_c3_clk),                                //                    c3.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.c4                 (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (3'b000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	vga_lt24_accelerometer_computer_jtag_uart_0 jtag_uart_0 (
		.clk            (altpll_0_c2_clk),                                             //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                             //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                                     //               irq.irq
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (8),
		.RESPONSE_FIFO_DEPTH (8),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge (
		.m0_clk           (altpll_0_c3_clk),                                             //   m0_clk.clk
		.m0_reset         (rst_controller_001_reset_out_reset),                          // m0_reset.reset
		.s0_clk           (altpll_0_c2_clk),                                             //   s0_clk.clk
		.s0_reset         (rst_controller_002_reset_out_reset),                          // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_m0_writedata),                       //         .writedata
		.m0_address       (mm_clock_crossing_bridge_m0_address),                         //         .address
		.m0_write         (mm_clock_crossing_bridge_m0_write),                           //         .write
		.m0_read          (mm_clock_crossing_bridge_m0_read),                            //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_m0_debugaccess)                      //         .debugaccess
	);

	vga_lt24_accelerometer_computer_new_sdram_controller_0 new_sdram_controller_0 (
		.clk            (altpll_0_c2_clk),                                           //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),                           // reset.reset_n
		.az_addr        (mm_interconnect_0_new_sdram_controller_0_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_new_sdram_controller_0_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_new_sdram_controller_0_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_new_sdram_controller_0_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_new_sdram_controller_0_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_new_sdram_controller_0_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                           //  wire.export
		.zs_ba          (sdram_wire_ba),                                             //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                          //      .export
		.zs_cke         (sdram_wire_cke),                                            //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                           //      .export
		.zs_dq          (sdram_wire_dq),                                             //      .export
		.zs_dqm         (sdram_wire_dqm),                                            //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                          //      .export
		.zs_we_n        (sdram_wire_we_n)                                            //      .export
	);

	vga_lt24_accelerometer_computer_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (altpll_0_c2_clk),                                            //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                            //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                         //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.d_burstcount                        (nios2_gen2_0_data_master_burstcount),                        //                          .burstcount
		.d_readdatavalid                     (nios2_gen2_0_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.i_burstcount                        (nios2_gen2_0_instruction_master_burstcount),                 //                          .burstcount
		.i_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	vga_lt24_accelerometer_computer_onchip_memory2_0 onchip_memory2_0 (
		.clk        (altpll_0_c2_clk),                                  //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_0_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_0_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_0_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_0_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_0_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_0_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_0_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),               //       .reset_req
		.freeze     (1'b0)                                              // (terminated)
	);

	vga_lt24_accelerometer_computer_sysid_qsys_0 sysid_qsys_0 (
		.clock    (altpll_0_c2_clk),                                       //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                       //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	vga_lt24_accelerometer_computer_timer_0 timer_0 (
		.clk        (altpll_0_c2_clk),                         //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver2_irq)                 //   irq.irq
	);

	vga_lt24_accelerometer_computer_timer_0 timer_1 (
		.clk        (altpll_0_c2_clk),                         //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_1_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_1_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_1_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_1_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_1_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver5_irq)                 //   irq.irq
	);

	vga_lt24_accelerometer_computer_touch_busy touch_busy (
		.clk      (altpll_0_c3_clk),                          //                 clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_1_touch_busy_s1_address),  //                  s1.address
		.readdata (mm_interconnect_1_touch_busy_s1_readdata), //                    .readdata
		.in_port  (touch_busy_external_connection_export)     // external_connection.export
	);

	vga_lt24_accelerometer_computer_touch_pen_irq_n touch_pen_irq_n (
		.clk        (altpll_0_c3_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_1_touch_pen_irq_n_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_touch_pen_irq_n_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_touch_pen_irq_n_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_touch_pen_irq_n_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_touch_pen_irq_n_s1_readdata),   //                    .readdata
		.in_port    (touch_pen_irq_n_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)                    //                 irq.irq
	);

	vga_lt24_accelerometer_computer_touch_spi touch_spi (
		.clk           (altpll_0_c3_clk),                                         //              clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),                     //            reset.reset_n
		.data_from_cpu (mm_interconnect_1_touch_spi_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_1_touch_spi_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_1_touch_spi_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_1_touch_spi_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_1_touch_spi_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_1_touch_spi_spi_control_port_write),     //                 .write_n
		.irq           (irq_synchronizer_001_receiver_irq),                       //              irq.irq
		.MISO          (spi_external_MISO),                                       //         external.export
		.MOSI          (spi_external_MOSI),                                       //                 .export
		.SCLK          (spi_external_SCLK),                                       //                 .export
		.SS_n          (spi_external_SS_n)                                        //                 .export
	);

	vga_lt24_accelerometer_computer_video_dual_clock_buffer_0 video_dual_clock_buffer_0 (
		.clk_stream_in            (altpll_0_c2_clk),                                                 //         clock_stream_in.clk
		.reset_stream_in          (rst_controller_reset_out_reset),                                  //         reset_stream_in.reset
		.clk_stream_out           (altpll_0_c0_clk),                                                 //        clock_stream_out.clk
		.reset_stream_out         (rst_controller_004_reset_out_reset),                              //        reset_stream_out.reset
		.stream_in_ready          (video_rgb_resampler_0_avalon_rgb_source_ready),                   //   avalon_dc_buffer_sink.ready
		.stream_in_startofpacket  (video_rgb_resampler_0_avalon_rgb_source_startofpacket),           //                        .startofpacket
		.stream_in_endofpacket    (video_rgb_resampler_0_avalon_rgb_source_endofpacket),             //                        .endofpacket
		.stream_in_valid          (video_rgb_resampler_0_avalon_rgb_source_valid),                   //                        .valid
		.stream_in_data           (video_rgb_resampler_0_avalon_rgb_source_data),                    //                        .data
		.stream_out_ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         // avalon_dc_buffer_source.ready
		.stream_out_startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                        .startofpacket
		.stream_out_endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                        .endofpacket
		.stream_out_valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                        .valid
		.stream_out_data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data)           //                        .data
	);

	vga_lt24_accelerometer_computer_video_pixel_buffer_dma_0 video_pixel_buffer_dma_0 (
		.clk                  (altpll_0_c2_clk),                                                            //                     clk.clk
		.reset                (rst_controller_reset_out_reset),                                             //                   reset.reset
		.master_readdatavalid (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),             // avalon_pixel_dma_master.readdatavalid
		.master_waitrequest   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),               //                        .waitrequest
		.master_address       (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),                   //                        .address
		.master_arbiterlock   (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                      //                        .lock
		.master_read          (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),                      //                        .read
		.master_readdata      (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                  //                        .readdata
		.slave_address        (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address),    //    avalon_control_slave.address
		.slave_byteenable     (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable), //                        .byteenable
		.slave_read           (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read),       //                        .read
		.slave_write          (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write),      //                        .write
		.slave_writedata      (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata),  //                        .writedata
		.slave_readdata       (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata),   //                        .readdata
		.stream_ready         (video_pixel_buffer_dma_0_avalon_pixel_source_ready),                         //     avalon_pixel_source.ready
		.stream_startofpacket (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),                 //                        .startofpacket
		.stream_endofpacket   (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),                   //                        .endofpacket
		.stream_valid         (video_pixel_buffer_dma_0_avalon_pixel_source_valid),                         //                        .valid
		.stream_data          (video_pixel_buffer_dma_0_avalon_pixel_source_data)                           //                        .data
	);

	vga_lt24_accelerometer_computer_video_rgb_resampler_0 video_rgb_resampler_0 (
		.clk                      (altpll_0_c2_clk),                                                   //               clk.clk
		.reset                    (rst_controller_reset_out_reset),                                    //             reset.reset
		.stream_in_startofpacket  (video_pixel_buffer_dma_0_avalon_pixel_source_startofpacket),        //   avalon_rgb_sink.startofpacket
		.stream_in_endofpacket    (video_pixel_buffer_dma_0_avalon_pixel_source_endofpacket),          //                  .endofpacket
		.stream_in_valid          (video_pixel_buffer_dma_0_avalon_pixel_source_valid),                //                  .valid
		.stream_in_ready          (video_pixel_buffer_dma_0_avalon_pixel_source_ready),                //                  .ready
		.stream_in_data           (video_pixel_buffer_dma_0_avalon_pixel_source_data),                 //                  .data
		.slave_read               (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read),     //  avalon_rgb_slave.read
		.slave_readdata           (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata), //                  .readdata
		.stream_out_ready         (video_rgb_resampler_0_avalon_rgb_source_ready),                     // avalon_rgb_source.ready
		.stream_out_startofpacket (video_rgb_resampler_0_avalon_rgb_source_startofpacket),             //                  .startofpacket
		.stream_out_endofpacket   (video_rgb_resampler_0_avalon_rgb_source_endofpacket),               //                  .endofpacket
		.stream_out_valid         (video_rgb_resampler_0_avalon_rgb_source_valid),                     //                  .valid
		.stream_out_data          (video_rgb_resampler_0_avalon_rgb_source_data)                       //                  .data
	);

	vga_lt24_accelerometer_computer_video_vga_controller_0 video_vga_controller_0 (
		.clk           (altpll_0_c0_clk),                                                 //                clk.clk
		.reset         (rst_controller_004_reset_out_reset),                              //              reset.reset
		.data          (video_dual_clock_buffer_0_avalon_dc_buffer_source_data),          //    avalon_vga_sink.data
		.startofpacket (video_dual_clock_buffer_0_avalon_dc_buffer_source_startofpacket), //                   .startofpacket
		.endofpacket   (video_dual_clock_buffer_0_avalon_dc_buffer_source_endofpacket),   //                   .endofpacket
		.valid         (video_dual_clock_buffer_0_avalon_dc_buffer_source_valid),         //                   .valid
		.ready         (video_dual_clock_buffer_0_avalon_dc_buffer_source_ready),         //                   .ready
		.VGA_CLK       (vga_output_CLK),                                                  // external_interface.export
		.VGA_HS        (vga_output_HS),                                                   //                   .export
		.VGA_VS        (vga_output_VS),                                                   //                   .export
		.VGA_BLANK     (vga_output_BLANK),                                                //                   .export
		.VGA_SYNC      (vga_output_SYNC),                                                 //                   .export
		.VGA_R         (vga_output_R),                                                    //                   .export
		.VGA_G         (vga_output_G),                                                    //                   .export
		.VGA_B         (vga_output_B)                                                     //                   .export
	);

	vga_lt24_accelerometer_computer_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c2_clk                                                   (altpll_0_c2_clk),                                                                     //                                             altpll_0_c2.clk
		.clk_0_clk_clk                                                     (clk_clk),                                                                             //                                               clk_0_clk.clk
		.altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset        (rst_controller_003_reset_out_reset),                                                  //    altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset_reset     (rst_controller_002_reset_out_reset),                                                  // mm_clock_crossing_bridge_s0_reset_reset_bridge_in_reset.reset
		.video_pixel_buffer_dma_0_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                                                      //    video_pixel_buffer_dma_0_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address                                  (nios2_gen2_0_data_master_address),                                                    //                                nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest                              (nios2_gen2_0_data_master_waitrequest),                                                //                                                        .waitrequest
		.nios2_gen2_0_data_master_burstcount                               (nios2_gen2_0_data_master_burstcount),                                                 //                                                        .burstcount
		.nios2_gen2_0_data_master_byteenable                               (nios2_gen2_0_data_master_byteenable),                                                 //                                                        .byteenable
		.nios2_gen2_0_data_master_read                                     (nios2_gen2_0_data_master_read),                                                       //                                                        .read
		.nios2_gen2_0_data_master_readdata                                 (nios2_gen2_0_data_master_readdata),                                                   //                                                        .readdata
		.nios2_gen2_0_data_master_readdatavalid                            (nios2_gen2_0_data_master_readdatavalid),                                              //                                                        .readdatavalid
		.nios2_gen2_0_data_master_write                                    (nios2_gen2_0_data_master_write),                                                      //                                                        .write
		.nios2_gen2_0_data_master_writedata                                (nios2_gen2_0_data_master_writedata),                                                  //                                                        .writedata
		.nios2_gen2_0_data_master_debugaccess                              (nios2_gen2_0_data_master_debugaccess),                                                //                                                        .debugaccess
		.nios2_gen2_0_instruction_master_address                           (nios2_gen2_0_instruction_master_address),                                             //                         nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                                         //                                                        .waitrequest
		.nios2_gen2_0_instruction_master_burstcount                        (nios2_gen2_0_instruction_master_burstcount),                                          //                                                        .burstcount
		.nios2_gen2_0_instruction_master_read                              (nios2_gen2_0_instruction_master_read),                                                //                                                        .read
		.nios2_gen2_0_instruction_master_readdata                          (nios2_gen2_0_instruction_master_readdata),                                            //                                                        .readdata
		.nios2_gen2_0_instruction_master_readdatavalid                     (nios2_gen2_0_instruction_master_readdatavalid),                                       //                                                        .readdatavalid
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_address          (video_pixel_buffer_dma_0_avalon_pixel_dma_master_address),                            //        video_pixel_buffer_dma_0_avalon_pixel_dma_master.address
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest      (video_pixel_buffer_dma_0_avalon_pixel_dma_master_waitrequest),                        //                                                        .waitrequest
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_read             (video_pixel_buffer_dma_0_avalon_pixel_dma_master_read),                               //                                                        .read
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata         (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdata),                           //                                                        .readdata
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid    (video_pixel_buffer_dma_0_avalon_pixel_dma_master_readdatavalid),                      //                                                        .readdatavalid
		.video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock             (video_pixel_buffer_dma_0_avalon_pixel_dma_master_lock),                               //                                                        .lock
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_address     (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_address),     //   accelerometer_spi_avalon_accelerometer_spi_mode_slave.address
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_write       (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_write),       //                                                        .write
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_read        (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_read),        //                                                        .read
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_readdata    (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_readdata),    //                                                        .readdata
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_writedata   (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_writedata),   //                                                        .writedata
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_byteenable  (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_byteenable),  //                                                        .byteenable
		.accelerometer_spi_avalon_accelerometer_spi_mode_slave_waitrequest (mm_interconnect_0_accelerometer_spi_avalon_accelerometer_spi_mode_slave_waitrequest), //                                                        .waitrequest
		.altpll_0_pll_slave_address                                        (mm_interconnect_0_altpll_0_pll_slave_address),                                        //                                      altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                                          (mm_interconnect_0_altpll_0_pll_slave_write),                                          //                                                        .write
		.altpll_0_pll_slave_read                                           (mm_interconnect_0_altpll_0_pll_slave_read),                                           //                                                        .read
		.altpll_0_pll_slave_readdata                                       (mm_interconnect_0_altpll_0_pll_slave_readdata),                                       //                                                        .readdata
		.altpll_0_pll_slave_writedata                                      (mm_interconnect_0_altpll_0_pll_slave_writedata),                                      //                                                        .writedata
		.HEX3_HEX0_s1_address                                              (mm_interconnect_0_hex3_hex0_s1_address),                                              //                                            HEX3_HEX0_s1.address
		.HEX3_HEX0_s1_write                                                (mm_interconnect_0_hex3_hex0_s1_write),                                                //                                                        .write
		.HEX3_HEX0_s1_readdata                                             (mm_interconnect_0_hex3_hex0_s1_readdata),                                             //                                                        .readdata
		.HEX3_HEX0_s1_writedata                                            (mm_interconnect_0_hex3_hex0_s1_writedata),                                            //                                                        .writedata
		.HEX3_HEX0_s1_chipselect                                           (mm_interconnect_0_hex3_hex0_s1_chipselect),                                           //                                                        .chipselect
		.HEX5_HEX4_s1_address                                              (mm_interconnect_0_hex5_hex4_s1_address),                                              //                                            HEX5_HEX4_s1.address
		.HEX5_HEX4_s1_write                                                (mm_interconnect_0_hex5_hex4_s1_write),                                                //                                                        .write
		.HEX5_HEX4_s1_readdata                                             (mm_interconnect_0_hex5_hex4_s1_readdata),                                             //                                                        .readdata
		.HEX5_HEX4_s1_writedata                                            (mm_interconnect_0_hex5_hex4_s1_writedata),                                            //                                                        .writedata
		.HEX5_HEX4_s1_chipselect                                           (mm_interconnect_0_hex5_hex4_s1_chipselect),                                           //                                                        .chipselect
		.jtag_uart_0_avalon_jtag_slave_address                             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),                             //                           jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write                               (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),                               //                                                        .write
		.jtag_uart_0_avalon_jtag_slave_read                                (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),                                //                                                        .read
		.jtag_uart_0_avalon_jtag_slave_readdata                            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),                            //                                                        .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata                           (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),                           //                                                        .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest                         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest),                         //                                                        .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect                          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),                          //                                                        .chipselect
		.KEY_s1_address                                                    (mm_interconnect_0_key_s1_address),                                                    //                                                  KEY_s1.address
		.KEY_s1_write                                                      (mm_interconnect_0_key_s1_write),                                                      //                                                        .write
		.KEY_s1_readdata                                                   (mm_interconnect_0_key_s1_readdata),                                                   //                                                        .readdata
		.KEY_s1_writedata                                                  (mm_interconnect_0_key_s1_writedata),                                                  //                                                        .writedata
		.KEY_s1_chipselect                                                 (mm_interconnect_0_key_s1_chipselect),                                                 //                                                        .chipselect
		.LEDS_s1_address                                                   (mm_interconnect_0_leds_s1_address),                                                   //                                                 LEDS_s1.address
		.LEDS_s1_write                                                     (mm_interconnect_0_leds_s1_write),                                                     //                                                        .write
		.LEDS_s1_readdata                                                  (mm_interconnect_0_leds_s1_readdata),                                                  //                                                        .readdata
		.LEDS_s1_writedata                                                 (mm_interconnect_0_leds_s1_writedata),                                                 //                                                        .writedata
		.LEDS_s1_chipselect                                                (mm_interconnect_0_leds_s1_chipselect),                                                //                                                        .chipselect
		.mm_clock_crossing_bridge_s0_address                               (mm_interconnect_0_mm_clock_crossing_bridge_s0_address),                               //                             mm_clock_crossing_bridge_s0.address
		.mm_clock_crossing_bridge_s0_write                                 (mm_interconnect_0_mm_clock_crossing_bridge_s0_write),                                 //                                                        .write
		.mm_clock_crossing_bridge_s0_read                                  (mm_interconnect_0_mm_clock_crossing_bridge_s0_read),                                  //                                                        .read
		.mm_clock_crossing_bridge_s0_readdata                              (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdata),                              //                                                        .readdata
		.mm_clock_crossing_bridge_s0_writedata                             (mm_interconnect_0_mm_clock_crossing_bridge_s0_writedata),                             //                                                        .writedata
		.mm_clock_crossing_bridge_s0_burstcount                            (mm_interconnect_0_mm_clock_crossing_bridge_s0_burstcount),                            //                                                        .burstcount
		.mm_clock_crossing_bridge_s0_byteenable                            (mm_interconnect_0_mm_clock_crossing_bridge_s0_byteenable),                            //                                                        .byteenable
		.mm_clock_crossing_bridge_s0_readdatavalid                         (mm_interconnect_0_mm_clock_crossing_bridge_s0_readdatavalid),                         //                                                        .readdatavalid
		.mm_clock_crossing_bridge_s0_waitrequest                           (mm_interconnect_0_mm_clock_crossing_bridge_s0_waitrequest),                           //                                                        .waitrequest
		.mm_clock_crossing_bridge_s0_debugaccess                           (mm_interconnect_0_mm_clock_crossing_bridge_s0_debugaccess),                           //                                                        .debugaccess
		.new_sdram_controller_0_s1_address                                 (mm_interconnect_0_new_sdram_controller_0_s1_address),                                 //                               new_sdram_controller_0_s1.address
		.new_sdram_controller_0_s1_write                                   (mm_interconnect_0_new_sdram_controller_0_s1_write),                                   //                                                        .write
		.new_sdram_controller_0_s1_read                                    (mm_interconnect_0_new_sdram_controller_0_s1_read),                                    //                                                        .read
		.new_sdram_controller_0_s1_readdata                                (mm_interconnect_0_new_sdram_controller_0_s1_readdata),                                //                                                        .readdata
		.new_sdram_controller_0_s1_writedata                               (mm_interconnect_0_new_sdram_controller_0_s1_writedata),                               //                                                        .writedata
		.new_sdram_controller_0_s1_byteenable                              (mm_interconnect_0_new_sdram_controller_0_s1_byteenable),                              //                                                        .byteenable
		.new_sdram_controller_0_s1_readdatavalid                           (mm_interconnect_0_new_sdram_controller_0_s1_readdatavalid),                           //                                                        .readdatavalid
		.new_sdram_controller_0_s1_waitrequest                             (mm_interconnect_0_new_sdram_controller_0_s1_waitrequest),                             //                                                        .waitrequest
		.new_sdram_controller_0_s1_chipselect                              (mm_interconnect_0_new_sdram_controller_0_s1_chipselect),                              //                                                        .chipselect
		.nios2_gen2_0_debug_mem_slave_address                              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),                              //                            nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write                                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),                                //                                                        .write
		.nios2_gen2_0_debug_mem_slave_read                                 (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),                                 //                                                        .read
		.nios2_gen2_0_debug_mem_slave_readdata                             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),                             //                                                        .readdata
		.nios2_gen2_0_debug_mem_slave_writedata                            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),                            //                                                        .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable                           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),                           //                                                        .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),                          //                                                        .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess                          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),                          //                                                        .debugaccess
		.onchip_memory2_0_s1_address                                       (mm_interconnect_0_onchip_memory2_0_s1_address),                                       //                                     onchip_memory2_0_s1.address
		.onchip_memory2_0_s1_write                                         (mm_interconnect_0_onchip_memory2_0_s1_write),                                         //                                                        .write
		.onchip_memory2_0_s1_readdata                                      (mm_interconnect_0_onchip_memory2_0_s1_readdata),                                      //                                                        .readdata
		.onchip_memory2_0_s1_writedata                                     (mm_interconnect_0_onchip_memory2_0_s1_writedata),                                     //                                                        .writedata
		.onchip_memory2_0_s1_byteenable                                    (mm_interconnect_0_onchip_memory2_0_s1_byteenable),                                    //                                                        .byteenable
		.onchip_memory2_0_s1_chipselect                                    (mm_interconnect_0_onchip_memory2_0_s1_chipselect),                                    //                                                        .chipselect
		.onchip_memory2_0_s1_clken                                         (mm_interconnect_0_onchip_memory2_0_s1_clken),                                         //                                                        .clken
		.SLIDERS_s1_address                                                (mm_interconnect_0_sliders_s1_address),                                                //                                              SLIDERS_s1.address
		.SLIDERS_s1_readdata                                               (mm_interconnect_0_sliders_s1_readdata),                                               //                                                        .readdata
		.sysid_qsys_0_control_slave_address                                (mm_interconnect_0_sysid_qsys_0_control_slave_address),                                //                              sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata                               (mm_interconnect_0_sysid_qsys_0_control_slave_readdata),                               //                                                        .readdata
		.timer_0_s1_address                                                (mm_interconnect_0_timer_0_s1_address),                                                //                                              timer_0_s1.address
		.timer_0_s1_write                                                  (mm_interconnect_0_timer_0_s1_write),                                                  //                                                        .write
		.timer_0_s1_readdata                                               (mm_interconnect_0_timer_0_s1_readdata),                                               //                                                        .readdata
		.timer_0_s1_writedata                                              (mm_interconnect_0_timer_0_s1_writedata),                                              //                                                        .writedata
		.timer_0_s1_chipselect                                             (mm_interconnect_0_timer_0_s1_chipselect),                                             //                                                        .chipselect
		.timer_1_s1_address                                                (mm_interconnect_0_timer_1_s1_address),                                                //                                              timer_1_s1.address
		.timer_1_s1_write                                                  (mm_interconnect_0_timer_1_s1_write),                                                  //                                                        .write
		.timer_1_s1_readdata                                               (mm_interconnect_0_timer_1_s1_readdata),                                               //                                                        .readdata
		.timer_1_s1_writedata                                              (mm_interconnect_0_timer_1_s1_writedata),                                              //                                                        .writedata
		.timer_1_s1_chipselect                                             (mm_interconnect_0_timer_1_s1_chipselect),                                             //                                                        .chipselect
		.video_pixel_buffer_dma_0_avalon_control_slave_address             (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_address),             //           video_pixel_buffer_dma_0_avalon_control_slave.address
		.video_pixel_buffer_dma_0_avalon_control_slave_write               (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_write),               //                                                        .write
		.video_pixel_buffer_dma_0_avalon_control_slave_read                (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_read),                //                                                        .read
		.video_pixel_buffer_dma_0_avalon_control_slave_readdata            (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_readdata),            //                                                        .readdata
		.video_pixel_buffer_dma_0_avalon_control_slave_writedata           (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_writedata),           //                                                        .writedata
		.video_pixel_buffer_dma_0_avalon_control_slave_byteenable          (mm_interconnect_0_video_pixel_buffer_dma_0_avalon_control_slave_byteenable),          //                                                        .byteenable
		.video_rgb_resampler_0_avalon_rgb_slave_read                       (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_read),                       //                  video_rgb_resampler_0_avalon_rgb_slave.read
		.video_rgb_resampler_0_avalon_rgb_slave_readdata                   (mm_interconnect_0_video_rgb_resampler_0_avalon_rgb_slave_readdata)                    //                                                        .readdata
	);

	vga_lt24_accelerometer_computer_mm_interconnect_1 mm_interconnect_1 (
		.altpll_0_c2_clk                                               (altpll_0_c2_clk),                                             //                                             altpll_0_c2.clk
		.altpll_0_c3_clk                                               (altpll_0_c3_clk),                                             //                                             altpll_0_c3.clk
		.LT24_Controller_reset_reset_bridge_in_reset_reset             (rst_controller_002_reset_out_reset),                          //             LT24_Controller_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // mm_clock_crossing_bridge_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_m0_address                           (mm_clock_crossing_bridge_m0_address),                         //                             mm_clock_crossing_bridge_m0.address
		.mm_clock_crossing_bridge_m0_waitrequest                       (mm_clock_crossing_bridge_m0_waitrequest),                     //                                                        .waitrequest
		.mm_clock_crossing_bridge_m0_burstcount                        (mm_clock_crossing_bridge_m0_burstcount),                      //                                                        .burstcount
		.mm_clock_crossing_bridge_m0_byteenable                        (mm_clock_crossing_bridge_m0_byteenable),                      //                                                        .byteenable
		.mm_clock_crossing_bridge_m0_read                              (mm_clock_crossing_bridge_m0_read),                            //                                                        .read
		.mm_clock_crossing_bridge_m0_readdata                          (mm_clock_crossing_bridge_m0_readdata),                        //                                                        .readdata
		.mm_clock_crossing_bridge_m0_readdatavalid                     (mm_clock_crossing_bridge_m0_readdatavalid),                   //                                                        .readdatavalid
		.mm_clock_crossing_bridge_m0_write                             (mm_clock_crossing_bridge_m0_write),                           //                                                        .write
		.mm_clock_crossing_bridge_m0_writedata                         (mm_clock_crossing_bridge_m0_writedata),                       //                                                        .writedata
		.mm_clock_crossing_bridge_m0_debugaccess                       (mm_clock_crossing_bridge_m0_debugaccess),                     //                                                        .debugaccess
		.LCD_RESET_N_s1_address                                        (mm_interconnect_1_lcd_reset_n_s1_address),                    //                                          LCD_RESET_N_s1.address
		.LCD_RESET_N_s1_write                                          (mm_interconnect_1_lcd_reset_n_s1_write),                      //                                                        .write
		.LCD_RESET_N_s1_readdata                                       (mm_interconnect_1_lcd_reset_n_s1_readdata),                   //                                                        .readdata
		.LCD_RESET_N_s1_writedata                                      (mm_interconnect_1_lcd_reset_n_s1_writedata),                  //                                                        .writedata
		.LCD_RESET_N_s1_chipselect                                     (mm_interconnect_1_lcd_reset_n_s1_chipselect),                 //                                                        .chipselect
		.LT24_Controller_avalon_slave_0_address                        (mm_interconnect_1_lt24_controller_avalon_slave_0_address),    //                          LT24_Controller_avalon_slave_0.address
		.LT24_Controller_avalon_slave_0_write                          (mm_interconnect_1_lt24_controller_avalon_slave_0_write),      //                                                        .write
		.LT24_Controller_avalon_slave_0_writedata                      (mm_interconnect_1_lt24_controller_avalon_slave_0_writedata),  //                                                        .writedata
		.LT24_Controller_avalon_slave_0_chipselect                     (mm_interconnect_1_lt24_controller_avalon_slave_0_chipselect), //                                                        .chipselect
		.touch_busy_s1_address                                         (mm_interconnect_1_touch_busy_s1_address),                     //                                           touch_busy_s1.address
		.touch_busy_s1_readdata                                        (mm_interconnect_1_touch_busy_s1_readdata),                    //                                                        .readdata
		.touch_pen_irq_n_s1_address                                    (mm_interconnect_1_touch_pen_irq_n_s1_address),                //                                      touch_pen_irq_n_s1.address
		.touch_pen_irq_n_s1_write                                      (mm_interconnect_1_touch_pen_irq_n_s1_write),                  //                                                        .write
		.touch_pen_irq_n_s1_readdata                                   (mm_interconnect_1_touch_pen_irq_n_s1_readdata),               //                                                        .readdata
		.touch_pen_irq_n_s1_writedata                                  (mm_interconnect_1_touch_pen_irq_n_s1_writedata),              //                                                        .writedata
		.touch_pen_irq_n_s1_chipselect                                 (mm_interconnect_1_touch_pen_irq_n_s1_chipselect),             //                                                        .chipselect
		.touch_spi_spi_control_port_address                            (mm_interconnect_1_touch_spi_spi_control_port_address),        //                              touch_spi_spi_control_port.address
		.touch_spi_spi_control_port_write                              (mm_interconnect_1_touch_spi_spi_control_port_write),          //                                                        .write
		.touch_spi_spi_control_port_read                               (mm_interconnect_1_touch_spi_spi_control_port_read),           //                                                        .read
		.touch_spi_spi_control_port_readdata                           (mm_interconnect_1_touch_spi_spi_control_port_readdata),       //                                                        .readdata
		.touch_spi_spi_control_port_writedata                          (mm_interconnect_1_touch_spi_spi_control_port_writedata),      //                                                        .writedata
		.touch_spi_spi_control_port_chipselect                         (mm_interconnect_1_touch_spi_spi_control_port_chipselect)      //                                                        .chipselect
	);

	vga_lt24_accelerometer_computer_irq_mapper irq_mapper (
		.clk           (altpll_0_c2_clk),                //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),       // receiver5.irq
		.sender_irq    (nios2_gen2_0_irq_irq)            //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (altpll_0_c3_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c2_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (altpll_0_c3_clk),                    //       receiver_clk.clk
		.sender_clk     (altpll_0_c2_clk),                    //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_0_c2_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req),     //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_0_c3_clk),                    //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (altpll_0_c2_clk),                    //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (altpll_0_c0_clk),                        //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),     // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
